entity addpc is 
pc_cu : in std_logic_vector (31 downto 0);
pc_ne: out std_logic_vector(31 downto 0);
end addpc;

architecture dtflow 
